let gmbs_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[gmbs]
let gm_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[gm]
let gds_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[gds]
let vdsat_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[vdsat]
let vth_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[vth]
let id_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[id]
let ibd_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[ibd]
let ibs_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[ibs]
let gbd_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[gbd]
let gbs_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[gbs]
let isub_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[isub]
let igidl_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[igidl]
let igisl_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[igisl]
let igs_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[igs]
let igd_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[igd]
let igb_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[igb]
let igcs_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[igcs]
let vbs_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[vbs]
let vgs_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[vgs]
let vds_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[vds]
let cgg_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[cgg]
let cgs_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[cgs]
let cgd_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[cgd]
let cbg_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[cbg]
let cbd_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[cbd]
let cbs_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[cbs]
let cdg_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[cdg]
let cdd_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[cdd]
let cds_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[cds]
let csg_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[csg]
let csd_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[csd]
let css_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[css]
let cgb_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[cgb]
let cdb_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[cdb]
let csb_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[csb]
let cbb_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[cbb]
let capbd_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[capbd]
let capbs_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[capbs]
let qg_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[qg]
let qb_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[qb]
let qs_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[qs]
let qinv_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[qinv]
let qdef_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[qdef]
let gcrg_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[gcrg]
let gtau_M1=@m.x1.x1.XM1.msky130_fd_pr__nfet_g5v0d10v5[gtau]

let gmbs_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[gmbs]
let gm_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[gm]
let gds_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[gds]
let vdsat_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[vdsat]
let vth_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[vth]
let id_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[id]
let ibd_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[ibd]
let ibs_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[ibs]
let gbd_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[gbd]
let gbs_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[gbs]
let isub_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[isub]
let igidl_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[igidl]
let igisl_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[igisl]
let igs_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[igs]
let igd_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[igd]
let igb_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[igb]
let igcs_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[igcs]
let vbs_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[vbs]
let vgs_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[vgs]
let vds_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[vds]
let cgg_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[cgg]
let cgs_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[cgs]
let cgd_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[cgd]
let cbg_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[cbg]
let cbd_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[cbd]
let cbs_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[cbs]
let cdg_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[cdg]
let cdd_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[cdd]
let cds_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[cds]
let csg_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[csg]
let csd_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[csd]
let css_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[css]
let cgb_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[cgb]
let cdb_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[cdb]
let csb_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[csb]
let cbb_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[cbb]
let capbd_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[capbd]
let capbs_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[capbs]
let qg_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[qg]
let qb_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[qb]
let qs_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[qs]
let qinv_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[qinv]
let qdef_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[qdef]
let gcrg_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[gcrg]
let gtau_M2=@m.x1.x1.XM2.msky130_fd_pr__nfet_g5v0d10v5[gtau]

let gmbs_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[gmbs]
let gm_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[gm]
let gds_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[gds]
let vdsat_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[vdsat]
let vth_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[vth]
let id_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[id]
let ibd_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[ibd]
let ibs_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[ibs]
let gbd_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[gbd]
let gbs_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[gbs]
let isub_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[isub]
let igidl_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[igidl]
let igisl_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[igisl]
let igs_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[igs]
let igd_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[igd]
let igb_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[igb]
let igcs_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[igcs]
let vbs_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[vbs]
let vgs_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[vgs]
let vds_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[vds]
let cgg_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[cgg]
let cgs_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[cgs]
let cgd_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[cgd]
let cbg_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[cbg]
let cbd_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[cbd]
let cbs_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[cbs]
let cdg_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[cdg]
let cdd_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[cdd]
let cds_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[cds]
let csg_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[csg]
let csd_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[csd]
let css_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[css]
let cgb_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[cgb]
let cdb_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[cdb]
let csb_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[csb]
let cbb_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[cbb]
let capbd_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[capbd]
let capbs_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[capbs]
let qg_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[qg]
let qb_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[qb]
let qs_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[qs]
let qinv_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[qinv]
let qdef_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[qdef]
let gcrg_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[gcrg]
let gtau_M3=@m.x1.x1.XM3.msky130_fd_pr__pfet_g5v0d10v5[gtau]

let gmbs_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[gmbs]
let gm_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[gm]
let gds_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[gds]
let vdsat_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[vdsat]
let vth_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[vth]
let id_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[id]
let ibd_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[ibd]
let ibs_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[ibs]
let gbd_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[gbd]
let gbs_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[gbs]
let isub_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[isub]
let igidl_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[igidl]
let igisl_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[igisl]
let igs_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[igs]
let igd_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[igd]
let igb_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[igb]
let igcs_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[igcs]
let vbs_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[vbs]
let vgs_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[vgs]
let vds_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[vds]
let cgg_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[cgg]
let cgs_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[cgs]
let cgd_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[cgd]
let cbg_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[cbg]
let cbd_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[cbd]
let cbs_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[cbs]
let cdg_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[cdg]
let cdd_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[cdd]
let cds_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[cds]
let csg_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[csg]
let csd_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[csd]
let css_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[css]
let cgb_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[cgb]
let cdb_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[cdb]
let csb_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[csb]
let cbb_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[cbb]
let capbd_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[capbd]
let capbs_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[capbs]
let qg_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[qg]
let qb_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[qb]
let qs_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[qs]
let qinv_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[qinv]
let qdef_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[qdef]
let gcrg_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[gcrg]
let gtau_M4=@m.x1.x1.XM4.msky130_fd_pr__pfet_g5v0d10v5[gtau]

let gmbs_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[gmbs]
let gm_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[gm]
let gds_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[gds]
let vdsat_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[vdsat]
let vth_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[vth]
let id_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[id]
let ibd_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[ibd]
let ibs_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[ibs]
let gbd_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[gbd]
let gbs_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[gbs]
let isub_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[isub]
let igidl_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[igidl]
let igisl_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[igisl]
let igs_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[igs]
let igd_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[igd]
let igb_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[igb]
let igcs_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[igcs]
let vbs_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[vbs]
let vgs_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[vgs]
let vds_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[vds]
let cgg_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[cgg]
let cgs_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[cgs]
let cgd_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[cgd]
let cbg_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[cbg]
let cbd_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[cbd]
let cbs_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[cbs]
let cdg_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[cdg]
let cdd_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[cdd]
let cds_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[cds]
let csg_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[csg]
let csd_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[csd]
let css_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[css]
let cgb_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[cgb]
let cdb_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[cdb]
let csb_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[csb]
let cbb_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[cbb]
let capbd_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[capbd]
let capbs_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[capbs]
let qg_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[qg]
let qb_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[qb]
let qs_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[qs]
let qinv_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[qinv]
let qdef_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[qdef]
let gcrg_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[gcrg]
let gtau_M5=@m.x1.x1.XM5.msky130_fd_pr__pfet_g5v0d10v5[gtau]

let gmbs_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[gmbs]
let gm_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[gm]
let gds_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[gds]
let vdsat_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[vdsat]
let vth_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[vth]
let id_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[id]
let ibd_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[ibd]
let ibs_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[ibs]
let gbd_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[gbd]
let gbs_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[gbs]
let isub_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[isub]
let igidl_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[igidl]
let igisl_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[igisl]
let igs_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[igs]
let igd_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[igd]
let igb_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[igb]
let igcs_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[igcs]
let vbs_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[vbs]
let vgs_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[vgs]
let vds_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[vds]
let cgg_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[cgg]
let cgs_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[cgs]
let cgd_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[cgd]
let cbg_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[cbg]
let cbd_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[cbd]
let cbs_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[cbs]
let cdg_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[cdg]
let cdd_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[cdd]
let cds_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[cds]
let csg_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[csg]
let csd_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[csd]
let css_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[css]
let cgb_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[cgb]
let cdb_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[cdb]
let csb_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[csb]
let cbb_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[cbb]
let capbd_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[capbd]
let capbs_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[capbs]
let qg_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[qg]
let qb_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[qb]
let qs_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[qs]
let qinv_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[qinv]
let qdef_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[qdef]
let gcrg_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[gcrg]
let gtau_M6=@m.x1.x1.XM6.msky130_fd_pr__pfet_g5v0d10v5[gtau]

let gmbs_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[gmbs]
let gm_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[gm]
let gds_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[gds]
let vdsat_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[vdsat]
let vth_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[vth]
let id_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[id]
let ibd_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[ibd]
let ibs_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[ibs]
let gbd_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[gbd]
let gbs_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[gbs]
let isub_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[isub]
let igidl_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[igidl]
let igisl_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[igisl]
let igs_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[igs]
let igd_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[igd]
let igb_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[igb]
let igcs_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[igcs]
let vbs_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[vbs]
let vgs_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[vgs]
let vds_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[vds]
let cgg_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[cgg]
let cgs_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[cgs]
let cgd_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[cgd]
let cbg_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[cbg]
let cbd_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[cbd]
let cbs_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[cbs]
let cdg_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[cdg]
let cdd_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[cdd]
let cds_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[cds]
let csg_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[csg]
let csd_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[csd]
let css_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[css]
let cgb_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[cgb]
let cdb_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[cdb]
let csb_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[csb]
let cbb_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[cbb]
let capbd_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[capbd]
let capbs_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[capbs]
let qg_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[qg]
let qb_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[qb]
let qs_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[qs]
let qinv_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[qinv]
let qdef_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[qdef]
let gcrg_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[gcrg]
let gtau_M7=@m.x1.x1.XM7.msky130_fd_pr__nfet_g5v0d10v5[gtau]

let gmbs_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[gmbs]
let gm_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[gm]
let gds_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[gds]
let vdsat_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[vdsat]
let vth_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[vth]
let id_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[id]
let ibd_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[ibd]
let ibs_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[ibs]
let gbd_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[gbd]
let gbs_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[gbs]
let isub_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[isub]
let igidl_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[igidl]
let igisl_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[igisl]
let igs_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[igs]
let igd_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[igd]
let igb_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[igb]
let igcs_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[igcs]
let vbs_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[vbs]
let vgs_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[vgs]
let vds_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[vds]
let cgg_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[cgg]
let cgs_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[cgs]
let cgd_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[cgd]
let cbg_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[cbg]
let cbd_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[cbd]
let cbs_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[cbs]
let cdg_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[cdg]
let cdd_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[cdd]
let cds_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[cds]
let csg_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[csg]
let csd_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[csd]
let css_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[css]
let cgb_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[cgb]
let cdb_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[cdb]
let csb_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[csb]
let cbb_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[cbb]
let capbd_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[capbd]
let capbs_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[capbs]
let qg_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[qg]
let qb_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[qb]
let qs_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[qs]
let qinv_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[qinv]
let qdef_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[qdef]
let gcrg_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[gcrg]
let gtau_M8=@m.x1.x1.XM8.msky130_fd_pr__nfet_g5v0d10v5[gtau]

let gmbs_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[gmbs]
let gm_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[gm]
let gds_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[gds]
let vdsat_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[vdsat]
let vth_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[vth]
let id_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[id]
let ibd_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[ibd]
let ibs_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[ibs]
let gbd_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[gbd]
let gbs_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[gbs]
let isub_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[isub]
let igidl_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[igidl]
let igisl_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[igisl]
let igs_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[igs]
let igd_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[igd]
let igb_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[igb]
let igcs_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[igcs]
let vbs_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[vbs]
let vgs_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[vgs]
let vds_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[vds]
let cgg_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[cgg]
let cgs_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[cgs]
let cgd_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[cgd]
let cbg_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[cbg]
let cbd_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[cbd]
let cbs_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[cbs]
let cdg_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[cdg]
let cdd_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[cdd]
let cds_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[cds]
let csg_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[csg]
let csd_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[csd]
let css_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[css]
let cgb_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[cgb]
let cdb_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[cdb]
let csb_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[csb]
let cbb_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[cbb]
let capbd_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[capbd]
let capbs_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[capbs]
let qg_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[qg]
let qb_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[qb]
let qs_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[qs]
let qinv_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[qinv]
let qdef_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[qdef]
let gcrg_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[gcrg]
let gtau_M9=@m.x1.x1.XM9.msky130_fd_pr__nfet_g5v0d10v5[gtau]

let gmbs_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[gmbs]
let gm_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[gm]
let gds_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[gds]
let vdsat_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[vdsat]
let vth_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[vth]
let id_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[id]
let ibd_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[ibd]
let ibs_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[ibs]
let gbd_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[gbd]
let gbs_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[gbs]
let isub_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[isub]
let igidl_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[igidl]
let igisl_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[igisl]
let igs_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[igs]
let igd_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[igd]
let igb_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[igb]
let igcs_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[igcs]
let vbs_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[vbs]
let vgs_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[vgs]
let vds_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[vds]
let cgg_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[cgg]
let cgs_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[cgs]
let cgd_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[cgd]
let cbg_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[cbg]
let cbd_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[cbd]
let cbs_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[cbs]
let cdg_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[cdg]
let cdd_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[cdd]
let cds_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[cds]
let csg_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[csg]
let csd_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[csd]
let css_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[css]
let cgb_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[cgb]
let cdb_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[cdb]
let csb_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[csb]
let cbb_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[cbb]
let capbd_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[capbd]
let capbs_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[capbs]
let qg_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[qg]
let qb_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[qb]
let qs_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[qs]
let qinv_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[qinv]
let qdef_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[qdef]
let gcrg_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[gcrg]
let gtau_M10=@m.x1.XM10.msky130_fd_pr__pfet_g5v0d10v5[gtau]

let dc_Vb1=@Vb1[dc]
let acmag_Vb1=@Vb1[acmag]
let acphase_Vb1=@Vb1[acphase]
let acreal_Vb1=@Vb1[acreal]
let acimag_Vb1=@Vb1[acimag]
let i_Vb1=@Vb1[i]
let p_Vb1=@Vb1[p]

let dc_Vb2=@Vb2[dc]
let acmag_Vb2=@Vb2[acmag]
let acphase_Vb2=@Vb2[acphase]
let acreal_Vb2=@Vb2[acreal]
let acimag_Vb2=@Vb2[acimag]
let i_Vb2=@Vb2[i]
let p_Vb2=@Vb2[p]

let capacitance_Cfb=@c.x1.XCfb.c1[capacitance]
let cap_Cfb=@c.x1.XCfb.c1[cap]
let c_Cfb=@c.x1.XCfb.c1[c]
let ic_Cfb=@c.x1.XCfb.c1[ic]
let temp_Cfb=@c.x1.XCfb.c1[temp]
let dtemp_Cfb=@c.x1.XCfb.c1[dtemp]
let w_Cfb=@c.x1.XCfb.c1[w]
let l_Cfb=@c.x1.XCfb.c1[l]
let m_Cfb=@c.x1.XCfb.c1[m]
let scale_Cfb=@c.x1.XCfb.c1[scale]
let i_Cfb=@c.x1.XCfb.c1[i]
let p_Cfb=@c.x1.XCfb.c1[p]
let sens_dc_Cfb=@c.x1.XCfb.c1[sens_dc]
let sens_real_Cfb=@c.x1.XCfb.c1[sens_real]
let sens_imag_Cfb=@c.x1.XCfb.c1[sens_imag]
let sens_mag_Cfb=@c.x1.XCfb.c1[sens_mag]
let sens_ph_Cfb=@c.x1.XCfb.c1[sens_ph]
let sens_cplx_Cfb=@c.x1.XCfb.c1[sens_cplx]

let capacitance_CL=@c.XCL.c1[capacitance]
let cap_CL=@c.XCL.c1[cap]
let c_CL=@c.XCL.c1[c]
let ic_CL=@c.XCL.c1[ic]
let temp_CL=@c.XCL.c1[temp]
let dtemp_CL=@c.XCL.c1[dtemp]
let w_CL=@c.XCL.c1[w]
let l_CL=@c.XCL.c1[l]
let m_CL=@c.XCL.c1[m]
let scale_CL=@c.XCL.c1[scale]
let i_CL=@c.XCL.c1[i]
let p_CL=@c.XCL.c1[p]
let sens_dc_CL=@c.XCL.c1[sens_dc]
let sens_real_CL=@c.XCL.c1[sens_real]
let sens_imag_CL=@c.XCL.c1[sens_imag]
let sens_mag_CL=@c.XCL.c1[sens_mag]
let sens_ph_CL=@c.XCL.c1[sens_ph]
let sens_cplx_CL=@c.XCL.c1[sens_cplx]

write ldo_folded_cascode_tb_op gmbs_M1 gm_M1 gds_M1 vdsat_M1 vth_M1 id_M1 ibd_M1 ibs_M1 gbd_M1 gbs_M1 isub_M1 igidl_M1 igisl_M1 igs_M1 igd_M1 igb_M1 igcs_M1 vbs_M1 vgs_M1 vds_M1 cgg_M1 cgs_M1 cgd_M1 cbg_M1 cbd_M1 cbs_M1 cdg_M1 cdd_M1 cds_M1 csg_M1 csd_M1 css_M1 cgb_M1 cdb_M1 csb_M1 cbb_M1 capbd_M1 capbs_M1 qg_M1 qb_M1 qs_M1 qinv_M1 qdef_M1 gcrg_M1 gtau_M1 gmbs_M2 gm_M2 gds_M2 vdsat_M2 vth_M2 id_M2 ibd_M2 ibs_M2 gbd_M2 gbs_M2 isub_M2 igidl_M2 igisl_M2 igs_M2 igd_M2 igb_M2 igcs_M2 vbs_M2 vgs_M2 vds_M2 cgg_M2 cgs_M2 cgd_M2 cbg_M2 cbd_M2 cbs_M2 cdg_M2 cdd_M2 cds_M2 csg_M2 csd_M2 css_M2 cgb_M2 cdb_M2 csb_M2 cbb_M2 capbd_M2 capbs_M2 qg_M2 qb_M2 qs_M2 qinv_M2 qdef_M2 gcrg_M2 gtau_M2 gmbs_M3 gm_M3 gds_M3 vdsat_M3 vth_M3 id_M3 ibd_M3 ibs_M3 gbd_M3 gbs_M3 isub_M3 igidl_M3 igisl_M3 igs_M3 igd_M3 igb_M3 igcs_M3 vbs_M3 vgs_M3 vds_M3 cgg_M3 cgs_M3 cgd_M3 cbg_M3 cbd_M3 cbs_M3 cdg_M3 cdd_M3 cds_M3 csg_M3 csd_M3 css_M3 cgb_M3 cdb_M3 csb_M3 cbb_M3 capbd_M3 capbs_M3 qg_M3 qb_M3 qs_M3 qinv_M3 qdef_M3 gcrg_M3 gtau_M3 gmbs_M4 gm_M4 gds_M4 vdsat_M4 vth_M4 id_M4 ibd_M4 ibs_M4 gbd_M4 gbs_M4 isub_M4 igidl_M4 igisl_M4 igs_M4 igd_M4 igb_M4 igcs_M4 vbs_M4 vgs_M4 vds_M4 cgg_M4 cgs_M4 cgd_M4 cbg_M4 cbd_M4 cbs_M4 cdg_M4 cdd_M4 cds_M4 csg_M4 csd_M4 css_M4 cgb_M4 cdb_M4 csb_M4 cbb_M4 capbd_M4 capbs_M4 qg_M4 qb_M4 qs_M4 qinv_M4 qdef_M4 gcrg_M4 gtau_M4 gmbs_M5 gm_M5 gds_M5 vdsat_M5 vth_M5 id_M5 ibd_M5 ibs_M5 gbd_M5 gbs_M5 isub_M5 igidl_M5 igisl_M5 igs_M5 igd_M5 igb_M5 igcs_M5 vbs_M5 vgs_M5 vds_M5 cgg_M5 cgs_M5 cgd_M5 cbg_M5 cbd_M5 cbs_M5 cdg_M5 cdd_M5 cds_M5 csg_M5 csd_M5 css_M5 cgb_M5 cdb_M5 csb_M5 cbb_M5 capbd_M5 capbs_M5 qg_M5 qb_M5 qs_M5 qinv_M5 qdef_M5 gcrg_M5 gtau_M5 gmbs_M6 gm_M6 gds_M6 vdsat_M6 vth_M6 id_M6 ibd_M6 ibs_M6 gbd_M6 gbs_M6 isub_M6 igidl_M6 igisl_M6 igs_M6 igd_M6 igb_M6 igcs_M6 vbs_M6 vgs_M6 vds_M6 cgg_M6 cgs_M6 cgd_M6 cbg_M6 cbd_M6 cbs_M6 cdg_M6 cdd_M6 cds_M6 csg_M6 csd_M6 css_M6 cgb_M6 cdb_M6 csb_M6 cbb_M6 capbd_M6 capbs_M6 qg_M6 qb_M6 qs_M6 qinv_M6 qdef_M6 gcrg_M6 gtau_M6 gmbs_M7 gm_M7 gds_M7 vdsat_M7 vth_M7 id_M7 ibd_M7 ibs_M7 gbd_M7 gbs_M7 isub_M7 igidl_M7 igisl_M7 igs_M7 igd_M7 igb_M7 igcs_M7 vbs_M7 vgs_M7 vds_M7 cgg_M7 cgs_M7 cgd_M7 cbg_M7 cbd_M7 cbs_M7 cdg_M7 cdd_M7 cds_M7 csg_M7 csd_M7 css_M7 cgb_M7 cdb_M7 csb_M7 cbb_M7 capbd_M7 capbs_M7 qg_M7 qb_M7 qs_M7 qinv_M7 qdef_M7 gcrg_M7 gtau_M7 gmbs_M8 gm_M8 gds_M8 vdsat_M8 vth_M8 id_M8 ibd_M8 ibs_M8 gbd_M8 gbs_M8 isub_M8 igidl_M8 igisl_M8 igs_M8 igd_M8 igb_M8 igcs_M8 vbs_M8 vgs_M8 vds_M8 cgg_M8 cgs_M8 cgd_M8 cbg_M8 cbd_M8 cbs_M8 cdg_M8 cdd_M8 cds_M8 csg_M8 csd_M8 css_M8 cgb_M8 cdb_M8 csb_M8 cbb_M8 capbd_M8 capbs_M8 qg_M8 qb_M8 qs_M8 qinv_M8 qdef_M8 gcrg_M8 gtau_M8 gmbs_M9 gm_M9 gds_M9 vdsat_M9 vth_M9 id_M9 ibd_M9 ibs_M9 gbd_M9 gbs_M9 isub_M9 igidl_M9 igisl_M9 igs_M9 igd_M9 igb_M9 igcs_M9 vbs_M9 vgs_M9 vds_M9 cgg_M9 cgs_M9 cgd_M9 cbg_M9 cbd_M9 cbs_M9 cdg_M9 cdd_M9 cds_M9 csg_M9 csd_M9 css_M9 cgb_M9 cdb_M9 csb_M9 cbb_M9 capbd_M9 capbs_M9 qg_M9 qb_M9 qs_M9 qinv_M9 qdef_M9 gcrg_M9 gtau_M9 gmbs_M10 gm_M10 gds_M10 vdsat_M10 vth_M10 id_M10 ibd_M10 ibs_M10 gbd_M10 gbs_M10 isub_M10 igidl_M10 igisl_M10 igs_M10 igd_M10 igb_M10 igcs_M10 vbs_M10 vgs_M10 vds_M10 cgg_M10 cgs_M10 cgd_M10 cbg_M10 cbd_M10 cbs_M10 cdg_M10 cdd_M10 cds_M10 csg_M10 csd_M10 css_M10 cgb_M10 cdb_M10 csb_M10 cbb_M10 capbd_M10 capbs_M10 qg_M10 qb_M10 qs_M10 qinv_M10 qdef_M10 gcrg_M10 gtau_M10 dc_Vb1 acmag_Vb1 acphase_Vb1 acreal_Vb1 acimag_Vb1 i_Vb1 p_Vb1 dc_Vb2 acmag_Vb2 acphase_Vb2 acreal_Vb2 acimag_Vb2 i_Vb2 p_Vb2 capacitance_Cfb cap_Cfb c_Cfb ic_Cfb temp_Cfb dtemp_Cfb w_Cfb l_Cfb m_Cfb scale_Cfb i_Cfb p_Cfb sens_dc_Cfb sens_real_Cfb sens_imag_Cfb sens_mag_Cfb sens_ph_Cfb sens_cplx_Cfb capacitance_CL cap_CL c_CL ic_CL temp_CL dtemp_CL w_CL l_CL m_CL scale_CL i_CL p_CL sens_dc_CL sens_real_CL sens_imag_CL sens_mag_CL sens_ph_CL sens_cplx_CL 
