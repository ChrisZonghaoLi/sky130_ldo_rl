.param W_M1=42.118154872134696 L_M1=1.7111959807328843
.param W_M2=42.118154872134696 L_M2=1.7111959807328843
.param W_M3=51.286530610841616 L_M3=2.5157359362276224
.param W_M4=51.286530610841616 L_M4=2.5157359362276224
.param W_M5=29.075754347959045 L_M5=1.6114024596504857
.param W_M6=57.71043983361096 L_M6=4.794129763236112
.param W_M7=13.16 L_M7=2.469795719604986
.param Rfb=2595.4894470684503 Cfb=1.837914159484712e-12
.param Vcm=0.7723338312726121 Vb=0.854368816484408
