.param W_M1=9.8838329911232 L_M1=1.3656668551266193
.param W_M2=W_M1 L_M2=L_M1
.param W_M3=81.09635359048843 L_M3=0.5364916324615479
.param W_M4=W_M3 L_M4=L_M3
.param W_M5=98.06255593895912 L_M5=0.6183840781450272
.param W_pass=20.553942620754242 L_pass=0.5468462407588959 M_pass=363
.param Vb=0.9322240442037582
.param M_Rfb=1 M_Cfb=7
.param M_CL=257
.param Vdd=2
.param Vref=1.8
.param IL=10m
