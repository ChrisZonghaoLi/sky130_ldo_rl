.param W_M1=72.18756159865863 L_M1=1.2410688308174198
.param W_M2=W_M1 L_M2=L_M1
.param W_M3=48.46762592099787 L_M3=1.8307155787659843
.param W_M4=W_M3 L_M4=L_M3
.param W_M5=83.2947084710894 L_M5=0.636778255202531
.param W_M6=W_M5 L_M6=L_M5
.param W_M7=77.86820461631672 L_M7=1.2423521011039824
.param W_M8=W_M7 L_M8=L_M7
.param W_M9=10.760224447365026 L_M9=0.5374729271299059
.param W_pass=28.750624611702865 L_pass=0.5917695569993786 M_pass=1461
.param Vb1=1.3450932697084956
.param Vb2=0.9099120399342119
.param M_Rfb=7
.param M_Cfb=36
.param M_CL=140
.param Vdd=2
.param Vref=1.8
.param IL=10m

