.param W_M1=12.286908000707626 L_M1=1.7774289548397064
.param W_M2=W_M1 L_M2=L_M1
.param W_M3=36.89915242791176 L_M3=0.5515819191932678
.param W_M4=W_M3 L_M4=L_M3
.param W_M5=12.32991936802864 L_M5=0.502713143825531
.param W_M6=W_M5 L_M6=L_M5
.param W_M7=91.40523833036423 L_M7=1.717549979686737
.param W_M8=W_M7 L_M8=L_M7
.param W_M9=32.27177633345127 L_M9=0.557290107011795
.param W_pass=11.55021220445633 L_pass=0.5032543540000916 M_pass=275
.param Vb1=0.9951694101095199
.param Vb2=0.02523776888847351
.param M_Rfb=1
.param M_Cfb=9
.param M_CL=239
.param Vdd=2
.param Vref=1.8
.param IL=10m


